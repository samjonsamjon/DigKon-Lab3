LIBRARY ieee;
USE ieee.std_logic_1164.all;
--use ieee.std_logic_unsigned.all;
USE std.textio.all;
USE ieee.numeric_std.all;

ENTITY procBus IS
	PORT(	INSTRUCTION	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		DATA		: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		ACC		: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		EXTDATA		: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		OUTPUT		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		ERR		: OUT STD_LOGIC;
		instrSEL	: IN STD_LOGIC;
		dataSEL		: IN STD_LOGIC;
		accSEL		: IN STD_LOGIC;
		extdataSEL	: IN STD_LOGIC);
end procBus;




ARCHITECTURE behavorial OF procBus IS
SIGNAL SELEC : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL SELOR1 : STD_LOGIC;
SIGNAL SELOR2 : STD_LOGIC;
SIGNAL SELOR3 : STD_LOGIC;
SIGNAL SELOR4 : STD_LOGIC;
SIGNAL SELOR5 : STD_LOGIC;
SIGNAL SELOR6 : STD_LOGIC;

SIGNAL ELR : STD_LOGIC;

BEGIN
SELEC(0) <= instrSEL;
SELEC(1) <= dataSEL;
SELEC(2) <= accSEL;
SELEC(3) <= extdataSEL;

SELOR1 <=	(SELEC(0) AND SELEC(1));
SELOR2 <=	(SELEC(0) AND SELEC(2));
SELOR3 <=	(SELEC(0) AND SELEC(3));
SELOR4 <=	(SELEC(1) AND SELEC(2));
SELOR5 <=	(SELEC(1) AND SELEC(3));
SELOR6 <=	(SELEC(2) AND SELEC(3));

ELR <= SELOR1 OR SELOR2 OR SELOR3 OR SELOR4 OR SELOR5 OR SELOR6;

ERR <= '1' WHEN ELR = '1' ELSE '0';

OUTPUT <= 	EXTDATA	WHEN SELEC(3) = '1' ELSE
		ACC 	WHEN SELEC(2) = '1' ELSE
		DATA 	WHEN SELEC(1) = '1' ELSE
		INSTRUCTION WHEN SELEC(0) = '1' ELSE
		"00000000";
END behavorial;